`include "uvm_macros.svh"
import uvm_pkg::*;

`include "intf.sv"
`include "mem.sv"
`include "mem_txn.sv"
`include "mem_seq.sv"
`include "mem_sqr.sv"
`include "mem_drv.sv"
`include "mem_mon.sv"
`include "mem_agt.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "mem_test.sv"