interface intf (input bit clk,rst);
  logic [3:0] a,b;
  logic       c;
  logic [4:0] sum;
endinterface