`include "uvm_macros.svh"
import uvm_pkg::*;

`include "intf.sv"
`include "adder.sv"
`include "adder_txn.sv"
`include "adder_seq.sv"
`include "adder_sqr.sv"
`include "adder_drv.sv"
`include "adder_mon.sv"
`include "adder_agt.sv"
`include "adder_sbd.sv"
`include "adder_env.sv"
`include "adder_test.sv"