class mem_test extends uvm_test;
  `uvm_component_utils(mem_test)

  mem_seq seq;
  mem_env env;

  function new(string name="mem_test",uvm_component parent);
    super.new(name,parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    seq = mem_seq::type_id::create("seq");
    env = mem_env::type_id::create("env",this);
  endfunction

  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
      seq.start(env.agt.sqr);
    phase.drop_objection(this);
    phase.phase_done.set_drain_time(this,50);
  endtask
endclass